magic
tech gf180mcuD
magscale 1 10
timestamp 1750740011
<< error_p >>
rect -34 69 -23 115
rect -118 -23 -107 23
rect 50 -23 61 23
rect -34 -115 -23 -69
<< pwell >>
rect -282 -246 282 246
<< nmos >>
rect -28 -22 28 22
<< ndiff >>
rect -120 23 -48 36
rect -120 -23 -107 23
rect -61 22 -48 23
rect 48 23 120 36
rect 48 22 61 23
rect -61 -22 -28 22
rect 28 -22 61 22
rect -61 -23 -48 -22
rect -120 -36 -48 -23
rect 48 -23 61 -22
rect 107 -23 120 23
rect 48 -36 120 -23
<< ndiffc >>
rect -107 -23 -61 23
rect 61 -23 107 23
<< psubdiff >>
rect -258 150 258 222
rect -258 106 -186 150
rect -258 -106 -245 106
rect -199 -106 -186 106
rect 186 106 258 150
rect -258 -150 -186 -106
rect 186 -106 199 106
rect 245 -106 258 106
rect 186 -150 258 -106
rect -258 -222 258 -150
<< psubdiffcont >>
rect -245 -106 -199 106
rect 199 -106 245 106
<< polysilicon >>
rect -36 115 36 128
rect -36 69 -23 115
rect 23 69 36 115
rect -36 56 36 69
rect -28 22 28 56
rect -28 -56 28 -22
rect -36 -69 36 -56
rect -36 -115 -23 -69
rect 23 -115 36 -69
rect -36 -128 36 -115
<< polycontact >>
rect -23 69 23 115
rect -23 -115 23 -69
<< metal1 >>
rect -245 163 245 209
rect -245 106 -199 163
rect -34 69 -23 115
rect 23 69 34 115
rect 199 106 245 163
rect -118 -23 -107 23
rect -61 -23 -50 23
rect 50 -23 61 23
rect 107 -23 118 23
rect -245 -163 -199 -106
rect -34 -115 -23 -69
rect 23 -115 34 -69
rect 199 -163 245 -106
rect -245 -209 245 -163
<< properties >>
string FIXED_BBOX -222 -186 222 186
string gencell nfet_03v3
string library gf180mcu
string parameters w 0.22 l 0.28 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
