magic
tech gf180mcuD
magscale 1 10
timestamp 1750740011
<< error_p >>
rect -48 53 -37 99
rect -125 -66 -79 18
rect 79 -66 125 18
<< pwell >>
rect -162 -136 162 136
<< nmos >>
rect -50 -68 50 20
<< ndiff >>
rect -138 7 -50 20
rect -138 -55 -125 7
rect -79 -55 -50 7
rect -138 -68 -50 -55
rect 50 7 138 20
rect 50 -55 79 7
rect 125 -55 138 7
rect 50 -68 138 -55
<< ndiffc >>
rect -125 -55 -79 7
rect 79 -55 125 7
<< polysilicon >>
rect -50 99 50 112
rect -50 53 -37 99
rect 37 53 50 99
rect -50 20 50 53
rect -50 -112 50 -68
<< polycontact >>
rect -37 53 37 99
<< metal1 >>
rect -48 53 -37 99
rect 37 53 48 99
rect -125 7 -79 18
rect -125 -66 -79 -55
rect 79 7 125 18
rect 79 -66 125 -55
<< properties >>
string gencell nfet_03v3
string library gf180mcu
string parameters w 0.44 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
