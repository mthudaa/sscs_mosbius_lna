magic
tech gf180mcuD
magscale 1 10
timestamp 1750740011
<< nwell >>
rect -224 -196 224 196
<< pmos >>
rect -50 -66 50 66
<< pdiff >>
rect -138 53 -50 66
rect -138 -53 -125 53
rect -79 -53 -50 53
rect -138 -66 -50 -53
rect 50 53 138 66
rect 50 -53 79 53
rect 125 -53 138 53
rect 50 -66 138 -53
<< pdiffc >>
rect -125 -53 -79 53
rect 79 -53 125 53
<< polysilicon >>
rect -50 66 50 110
rect -50 -110 50 -66
<< metal1 >>
rect -125 53 -79 64
rect -125 -64 -79 -53
rect 79 53 125 64
rect 79 -64 125 -53
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 0.66 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
